module top ();
	wire _w2_ ;
	LUT0 name0 (
		_w2_
	);
	defparam name0.INIT = 1'h0;

endmodule